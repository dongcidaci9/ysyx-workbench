module ysyx_23060201_IFU(
	input [31:0] pc_in,
	output [31:0] pc_out,
	output [31:0] inst
);

	assign pc_out = pc_in;

endmodule
